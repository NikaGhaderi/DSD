library verilog;
use verilog.vl_types.all;
entity tcam_TB is
end tcam_TB;
