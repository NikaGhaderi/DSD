library verilog;
use verilog.vl_types.all;
entity tcam_TB2 is
end tcam_TB2;
