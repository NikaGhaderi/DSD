library verilog;
use verilog.vl_types.all;
entity tcam_TB3 is
end tcam_TB3;
